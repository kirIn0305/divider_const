/*================================================================================
| Project name
|---------------------------------------------------------------------------------
| Block name  : divider_5_22
| Version     : 0.0.0
| Description : 
|     - const unsigned value divider (if you want use signed, you should calculate abs)
|     - i1 / i2 = o1  (i2 = const value)
|     - convert calculation method from divider to multiplier
|     - reference LSI/FPGAの回路アーキテクチャ設計法 P289
|---------------------------------------------------------------------------------
| Created by kirIn : author's email address
\===============================================================================*/

module divider_5_22(i1, o1);

//================================================================================
// Constants
//================================================================================
    parameter  BWI1 = 5;
    parameter  BWI2 = 10;
    parameter  BWO1 = 5;
    parameter  CONST_MULTI = 'b0000101111;

//================================================================================
// Declare Input and Output Pins
//================================================================================
    input [BWI1-1:0] i1;
    output [BWO1-1:0] o1;

//================================================================================
// Declare Wires and Regs
//================================================================================
    wire [BWI2-1:0] i2;
    wire [BWI1+BWI2-1:0] o_tmp;

//================================================================================
// Divider (To tell the Truth -> Multipiler)
//================================================================================
    assign i2 = CONST_MULTI;
    assign o_tmp = i1 * i2;

    assign o1 = o_tmp[BWI1+BWI2-1 : BWI1+BWI2-5];

endmodule